version https://git-lfs.github.com/spec/v1
oid sha256:03257aef91d0c3f4b47d50cec4a5cd8a4fd17828e33e7cac360c35e0c06cfdcf
size 2160
