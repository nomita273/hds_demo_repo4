version https://git-lfs.github.com/spec/v1
oid sha256:3861720ec0e2005156ed7fb53937c10ecb843673446a5096ea99da7657e13e6b
size 2245
