version https://git-lfs.github.com/spec/v1
oid sha256:3386e0bb3d3f4da559b229e3770250991c2bb877f25a532e393d5b43f9785983
size 6542
