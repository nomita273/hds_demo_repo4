version https://git-lfs.github.com/spec/v1
oid sha256:cfcb324feb05905468487bce78b1b44f2b3434b6040fdb255f7236043178fae7
size 2697
