version https://git-lfs.github.com/spec/v1
oid sha256:6263d4db8bb432a422c7517db8c1e5a276d0565ad3ef03d7f42238e179c34889
size 3762
