version https://git-lfs.github.com/spec/v1
oid sha256:2641000312c9c7aea56ef5c3977393a463fda1bfcbf708bf2fcb3ab3a28d155a
size 13419
