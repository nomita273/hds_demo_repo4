version https://git-lfs.github.com/spec/v1
oid sha256:e0bdd0486ade21a64622a74f19e749d54086b2d631a86442cdd6bae970e53c7d
size 3406
