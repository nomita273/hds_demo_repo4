version https://git-lfs.github.com/spec/v1
oid sha256:3c016ab6c1b088d5f291e687aa039f07f98d36770b1531a988248f48094f10d3
size 2760
