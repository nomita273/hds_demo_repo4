version https://git-lfs.github.com/spec/v1
oid sha256:4c52163bd02abb49a7e7eb71d5cdcca294ecd5a6e30f3b2f06c4c6c6d4b868bc
size 6084
