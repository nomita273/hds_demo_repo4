version https://git-lfs.github.com/spec/v1
oid sha256:1d0f89e3151e999abb0efdaba2e71ce18ef692d3999076358c2dda6372b872f6
size 6739
