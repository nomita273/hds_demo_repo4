version https://git-lfs.github.com/spec/v1
oid sha256:645493c76ce342b5ccb822fd545d0ac20d4fdd271b385b2e03ff6524bdb6a3d9
size 10518
