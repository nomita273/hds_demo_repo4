version https://git-lfs.github.com/spec/v1
oid sha256:b0f420bb382ccb55bad921cfa22731afcc943a00fb20a40228ec3de824af6954
size 8077
